package test_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"

`include "uart_xtn.sv"
`include "uart_agent_config.sv"
`include "env_config.sv"
`include "uart_driver.sv"
`include "uart_monitor.sv"
`include "uart_sequencer.sv"
`include "uart_agent.sv"
`include "uart_agent_top.sv"
`include "uart_seq.sv"

`include "virtual_sequencer.sv"
`include "virtual_seq.sv"
`include "scoreboard.sv"

`include "tb.sv"


`include "vtest_lib.sv"
endpackage
